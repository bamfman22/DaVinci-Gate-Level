// Name: alu.v
// Module: ALU
// Input: OP1[32] - operand 1
//        OP2[32] - operand 2
//        OPRN[6] - operation code
// Output: OUT[32] - output result for the operation
//
// Notes: 32 bit combinatorial ALU
// 
// Supports the following functions
//	- Integer add (0x1), sub(0x2), mul(0x3)
//	- Integer shift_rigth (0x4), shift_left (0x5)
//	- Bitwise and (0x6), or (0x7), nor (0x8)
//  - set less than (0x9)
//
// Revision History:
//
// Version	Date		Who		email			note
//------------------------------------------------------------------------------------------
//  1.0     Sep 10, 2014	Kaushik Patra	kpatra@sjsu.edu		Initial creation
//------------------------------------------------------------------------------------------
//
`include "prj_definition.v"
module ALU(OUT, ZERO, OP1, OP2, OPRN);
// input list
input [`DATA_INDEX_LIMIT:0] OP1; // operand 1
input [`DATA_INDEX_LIMIT:0] OP2; // operand 2
input [`ALU_OPRN_INDEX_LIMIT:0] OPRN; // operation code

// output list
output [`DATA_INDEX_LIMIT:0] OUT; // result of the operation.
output ZERO;

// TBD
wire [31:0] addSubWire;
wire [31:0] shiftWire;
wire [31:0] mulWire;
wire [31:0] andWire;
wire [31:0] orWire;
wire [31:0] norWire;
wire [31:0] muxWire;
wire [31:0] hiWire, test;
wire inv, and1, sna;

NOR32_2x1 n(norWire, OP1, OP2);

OR32_2x1  o(orWire, OP1, OP2);

AND32_2x1 a(andWire, OP1, OP2);

not invInit(inv, OPRN[0]);
and and1Init(and1, OPRN[3], OPRN[0]); 
or snaInit(sna, inv, and1);

RC_ADD_SUB_32 addSub(addSubWire, hiWire[0], OP1, OP2, sna);
MULT32 mul(hiWire, mulWire, OP1, OP2);
SHIFT32 shift(shiftWire, OP1, OP2, inv);


MUX32_16x1 mux(muxWire, addSubWire, addSubWire, addSubWire,
 mulWire, shiftWire, shiftWire, andWire, orWire,
 norWire, addSubWire, addSubWire, addSubWire, addSubWire,
 addSubWire, addSubWire, addSubWire, OPRN[3:0]);

BUF32_2x1 b(OUT, muxWire);

genvar i;
generate
	for(i = 0; i <32; i = i+1)
	begin : or_loop
		if(i == 31) begin
			or r(ZERO, test[i -1], 1'b0);
		end else if (i == 0) begin
			or r2(test[i], 1'b0, muxWire[i]);
		end else begin
			or r1(test[i], test[i-1], muxWire[i]);
		end
	end
endgenerate


endmodule
