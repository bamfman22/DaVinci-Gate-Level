
`timescale 1ns/1ps
module a_mux_tb;
	reg operand1, operand2, control;

	wire result;

	MUX1_2x1 m1(result, operand1,
		operand2, control);
	initial begin
		#5 control=0; operand1=0; operand2=0;
		#5 control=0; operand1=1; operand2=0;
		#5 control=0; operand1=0; operand2=1;
		#5 control=0; operand1=1; operand2=1;
		#5 control=1; operand1=0; operand2=0;
		#5 control=1; operand1=1; operand2=0;
		#5 control=1; operand1=0; operand2=1;
		#5 control=1; operand1=1; operand2=1;
	end
endmodule




module a_mux32_2x1_tb;


reg [31:0] I0,I1;
reg S;

wire [31:0] Y;

MUX32_2x1 m(Y,I0, I1, S);


initial begin
	#5 I0=15; I1 =12; S = 0;
	#5 I0 = 15; I1 =12; S=1;
end

endmodule

module a_32mux_tb;

reg[31:0]  I0, I1, I2, I3, I4, I5, I6, I7,
     I8, I9, I10, I11, I12, I13, I14, I15,
     I16, I17, I18, I19, I20, I21, I22, I23,
     I24, I25, I26, I27, I28, I29, I30, I31;

reg [4:0] S;


wire [31:0] Y;

MUX32_32x1 m(Y, I0, I1, I2, I3, I4, I5, I6, I7,
                     I8, I9, I10, I11, I12, I13, I14, I15,
                     I16, I17, I18, I19, I20, I21, I22, I23,
                     I24, I25, I26, I27, I28, I29, I30, I31, S);

initial begin
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =0;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =1;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =2;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =3;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =4;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =5;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =6;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =7;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =8;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =10;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =11;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =12;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =13;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =14;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =15;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =16;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =17;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =18;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =19;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =20;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =21;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =22;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =23;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =24;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =25;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =26;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =27;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =28;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =29;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =30;
	#5 I0 =10; I1=11; I2 = 12; I3=13; I4=14; I5=15; I6=16; I7=17; I8=18; I9=19; I10=110; I11=111; I12=112; I13=113; I14=114; I15=115; I16=116; I17=117; I18=118; I19=119; I20=210; I21=211; I22=212; I23=213;I24=214; I25=215; I26=216; I27=217; I28=218; I29=219; I30=310; I31=311; S =31;


	

end


endmodule

